LIBRARY ieee;
use ieee.std_logic_1164.all;
--------------------------------------------------------------------------------------------------------------------------
PACKAGE my_data_types IS
        TYPE matrix IS ARRAY (NATURAL RANGE <>, NATURAL RANGE <>) OF STD_LOGIC;
END PACKAGE my_data_types;
--------------------------------------------------------------------------------------------------------------------------
 