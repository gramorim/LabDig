library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;


entity operacoes_campo_fd is
	generic( constant ratio 		: integer := 434;
				constant log2_ratio 	: integer := 9;
				constant tam_ascii : integer := 7;
				constant filename : string := "campo_inicial.mif");
    port (
        clock, reset: in std_logic;
        partida : in std_logic;                    	-- tx_serial
        we: in std_logic;                          	-- memoria_jogo_16x7
        conta, zera, carrega: in std_logic;        	-- contador_m_load
        endereco: in std_logic_vector(5 downto 0); 	-- contador_m_load
        dado, sel: in std_logic_vector(1 downto 0);   -- mux3x1_n
        fim, fim_linha: out std_logic;             	-- contador_m_load
        saida_serial, pronto : out std_logic;      	-- tx_serial
        db_q: out std_logic_vector(5 downto 0);
        db_dados: out std_logic_vector(tam_ascii-1 downto 0);
        verifica: out std_logic_vector(1 downto 0);
		  i_verifica : in std_logic;
		  editavel : in std_logic
    );
end operacoes_campo_fd;

architecture operacoes_campo_fd of operacoes_campo_fd is
    signal s_contagem: std_logic_vector(5 downto 0);
    signal s_dados, s_mux, s_entrada: std_logic_vector (tam_ascii-1 downto 0);
	 signal s_verifica : std_logic_vector(1 downto 0);
	 signal s_fim4, s_fim8 : STD_LOGIC;

    component tx_serial 
	generic( constant ratio 		: integer;
				constant log2_ratio 	: integer;
				constant tam_ascii : integer);
				
   port(	clock, reset, partida, paridade	: in  std_logic;
			dados_ascii								: in  std_logic_vector (tam_ascii-1 downto 0);
			saida_serial, pronto 				: out std_logic;
			db_tick									: out std_logic);
    end component;
    
    component memoria_jogo_64x7 
	generic(	constant tam_ascii : integer;
				constant filename : string);
   PORT (dado_entrada : IN  STD_LOGIC_VECTOR(tam_ascii-1 DOWNTO 0);
         dado_saida   : OUT STD_LOGIC_VECTOR(tam_ascii-1 DOWNTO 0);
         endereco     : IN  STD_LOGIC_VECTOR(5 DOWNTO 0);         
         we, ce       : IN  STD_LOGIC);
    end component;

    component contador_m_load
    generic (
        constant M: integer;  -- modulo do contador
        constant N: integer   -- numero de bits da saida
    );
    port (
        CLK, zera, conta, carrega: in STD_LOGIC;
        D: in STD_LOGIC_VECTOR (N-1 downto 0);
        Q: out STD_LOGIC_VECTOR (N-1 downto 0);
        fim: out STD_LOGIC );
    end component;
    
    component mux3x1_n
      generic (
           constant BITS: integer);
      port(D2, D1, D0 : in std_logic_vector (BITS-1 downto 0);
           SEL: in std_logic_vector (1 downto 0);
           MX_OUT : out std_logic_vector (BITS-1 downto 0));
    end component;

    component decoder
		generic(constant tam_ascii : integer);
    port(
        input: in std_logic_vector (tam_ascii-1 downto 0);
        output : out std_logic_vector(1 downto 0)
    );
  end component; 
  
	component registrador_n is
	  generic (constant N: integer := 7);
	  port (clock, clear, enable: in STD_LOGIC;
			  D: in STD_LOGIC_VECTOR(N-1 downto 0);
			  Q: out STD_LOGIC_VECTOR (N-1 downto 0));
	end component;

	signal s_fim_linha, s_fim_coluna4, s_fim_coluna8, s_fim_coluna : std_logic;
begin

    -- sinais reset e partida mapeados em botoes ativos em alto
    U1: tx_serial 
		generic map(ratio,log2_ratio,tam_ascii)
		port map (clock=>clock, reset=>reset, partida=>partida, paridade=>'0',
                            dados_ascii=>s_mux, saida_serial=>saida_serial, pronto=>pronto);
    U2: memoria_jogo_64x7 
		generic map(tam_ascii,filename)
		PORT map(s_entrada,
					s_dados,
					s_contagem,        
					we, not editavel);
	
    U3: contador_m_load generic map (M => 64, N => 6) port map (CLK=>clock, zera=>zera, conta=>conta, carrega=>carrega,
                                                           D=>endereco, q=>s_contagem, fim=>fim);
    
	 --versao 7 bits
	 -- mux da saida memoria
    U4: mux3x1_n generic map (BITS => 7) port map (D2 => "0001101", D1=> "0001010", D0=>s_dados, 
                                                   SEL=>sel, MX_OUT=>s_mux);

    -- mux da entrada da memoria
    U5: mux3x1_n generic map (BITS => 7) port map (D2 => "1011000", D1=> "1000001", D0=>"1011111", 
                                                   SEL=>dado, MX_OUT=>s_entrada);
    
	-- versão 8 bits
	-- U4: mux3x1_n generic map (BITS => 8) port map (D2 => "10001101", D1=> "10001010", D0=>s_dados, 
   --                                                SEL=>sel, MX_OUT=>s_mux);

    -- mux da entrada da memoria
    --U5: mux3x1_n generic map (BITS => 8) port map (D2 => "11011000", D1=> "11000001", D0=>"11011111", 
    --                                               SEL=>dado, MX_OUT=>s_entrada);
   		 
    U6: decoder 
		generic map(tam_ascii)
		port map (input => s_dados, output => s_verifica);
	 
	 
	REG : registrador_n
	  generic map(2)
	  port map(clock, '0', i_verifica,
			  s_verifica,
			  verifica);

    with s_contagem(2 downto 0) select
        s_fim8 <= '1' when "111", '0' when others;
	with s_contagem(1 downto 0) select
			s_fim4 <= '1' when "11", '0' when others;
	with tamanho_campo select
			s_FIM_LINHA <= s_fim4 when '0', s_fim8 when '1';
			
			fim_linha <= s_fim_linha;

	with s_contagem(5 downto 3) select
		s_fim_coluna8 <= '1' when "111", '0' when others;

	with s_contagem(4 downto 3) select
		s_fim_coluna4 <= '1' when "11", '0' when others;
		
	

	with tamanho_campo select
		s_fim_coluna <= s_fim_coluna4 when '0', s_fim_coluna8 when '1';
	
	fim <= s_fim_coluna and s_fim_linha;
		
		
-- depuracao
db_q <= s_contagem;
db_dados <= s_mux;
    
end operacoes_campo_fd;

